module df();

endmodule